-- A DUT entity is used to wrap your design so that we can combine it with testbench.
-- This example shows how you can do this for the OR Gate

library ieee;
use ieee.std_logic_1164.all;

entity DUT is
    port(input_vector: in std_logic_vector(1 downto 0);
       	output_vector: out std_logic_vector(1 downto 0));
end entity;

architecture DutWrap of DUT is
   component ClockDivider is
     port (
    clk_in  : in  std_logic;
    rst   : in  std_logic;
    clk_out : out std_logic
);

   end component;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: ClockDivider
			port map (
    clk_in => input_vector(1),
    rst => input_vector(0),
    clk_out => output_vector(0)
);

end DutWrap;